library verilog;
use verilog.vl_types.all;
entity trabFinal_vlg_vec_tst is
end trabFinal_vlg_vec_tst;
